package riscv_pkg;

import uvm_pkg::*;

`include "remuldefs.svh"
`include "riscv_transaction.sv"
`include "riscv_sequence.sv"
`include "riscv_sequencer.sv"
`include "riscv_driver.sv"
`include "riscv_scoreboard.sv"
`include "riscv_agent.sv"
`include "riscv_environment.sv"
`include "riscv_test.sv"
`include "remul.sv"
//`include "dut_file"
`include "dut38.svp"
endpackage
